`timescale 1ns / 1ps

/*
 * Author:		李扬名.
 * StartTime:	18/11/9
 * Software:	Xilins-ISE
 * Editor:		Sublime
 * FileName:	Instr_ROM.v
 * FileType:	source
 * LastModify:	18/11/9
 */

 
module test_Data_ROM(
    );


endmodule
